module UART_MODULE_TB;
  localparam  WORD_LENGHT = 8;
   // Input Ports
  reg clk = 0;
  reg reset = 1;
  reg send = 0;
  reg value=1;

  reg [7:0]numero = 8'b1101_1011;

  UART_MODULE   DUT(
  	//Input Ports.
  	.clk_low(clk), .clk_high(clk),
  	.reset(reset),
  	.Rx_in(value),
  	.pop(1'b0),
  	.output_fifo_value(8'b1010_1010),

  	//Output Ports.
  	.Tx_out(),
  	.v(),
  	.fifos_out(),
  	.start(),
  	.fifo_out_pop(),
  	.n()

  );

  /*********************************************************/
  initial // Clock generator
    begin
      forever #2 clk = !clk;
    end
  /*********************************************************/
  initial begin // reset generator
  	#0 reset = 1;
    #4 reset = 0;
  	#4 reset = 1;
  end

  initial
    begin
    #200
      //Start
      //---------------------------Comando 1------------------------------
      #4 value = 0;
         numero = 'hFE;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //L
      #40 value = 0;
         numero = 'h3;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //CMD
      #40 value = 0;
         numero = 'h01;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //N
      #40 value = 0;
         numero = 'h4;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //END
      #40 value = 0;
         numero = 'hEF;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;

      //---------------------------Comando 2------------------------------
      #100
      //Start
      #4 value = 0;
         numero = 'hFE;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //L
      #40 value = 0;
         numero = 'h01;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //CMD
      #40 value = 0;
         numero = 'h02;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
      //END
      #40 value = 0;
         numero = 'hEF;
      #4  value = numero[0];
      #4  value = numero[1];
      #4  value = numero[2];
      #4  value = numero[3];
      #4  value = numero[4];
      #4  value = numero[5];
      #4  value = numero[6];
      #4  value = numero[7];
      #4 value = ^numero;
      #4 value = 1;
    end

endmodule
